library verilog;
use verilog.vl_types.all;
entity AluControlTestBench is
end AluControlTestBench;
