module or_32_bit(input [31:0] A , input [31:0] B , output [31:0] OUT);

or OR1(OUT[0], A[0] , B[0]);
or OR2(OUT[1], A[1] , B[1]);
or OR3(OUT[2], A[2] , B[2]);
or OR4(OUT[3], A[3] , B[3]);
or OR5(OUT[4], A[4] , B[4]);
or OR6(OUT[5], A[5] , B[5]);
or OR7(OUT[6], A[6] , B[6]);
or OR8(OUT[7], A[7] , B[7]);
or OR9(OUT[8], A[8] , B[8]);
or OR10(OUT[9], A[9] , B[9]);
or OR11(OUT[10], A[10] , B[10]);
or OR12(OUT[11], A[11] , B[11]);
or OR13(OUT[12], A[12] , B[12]);
or OR14(OUT[13], A[13] , B[13]);
or OR15(OUT[14], A[14] , B[14]);
or OR16(OUT[15], A[15] , B[15]);
or OR17(OUT[16], A[16] , B[16]);
or OR18(OUT[17], A[17] , B[17]);
or OR19(OUT[18], A[18] , B[18]);
or OR20(OUT[19], A[19] , B[19]);
or OR21(OUT[20], A[20] , B[20]);
or OR22(OUT[21], A[21] , B[21]);
or OR23(OUT[22], A[22] , B[22]);
or OR24(OUT[23], A[23] , B[23]);
or OR25(OUT[24], A[24] , B[24]);
or OR26(OUT[25], A[25] , B[25]);
or OR27(OUT[26], A[26] , B[26]);
or OR28(OUT[27], A[27] , B[27]);
or OR29(OUT[28], A[28] , B[28]);
or OR30(OUT[29], A[29] , B[29]);
or OR31(OUT[30], A[30] , B[30]);
or OR32(OUT[31], A[31] , B[31]);



endmodule