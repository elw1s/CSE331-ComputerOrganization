library verilog;
use verilog.vl_types.all;
entity not_32_bit_testbench is
end not_32_bit_testbench;
