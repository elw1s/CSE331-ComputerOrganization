library verilog;
use verilog.vl_types.all;
entity DataMemoryTestBench is
end DataMemoryTestBench;
