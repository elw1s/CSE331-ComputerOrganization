module and_32_bit(input [31:0] A , input [31:0] B , output [31:0] OUT);

and and1(OUT[0], A[0] , B[0]);
and and2(OUT[1], A[1] , B[1]);
and and3(OUT[2], A[2] , B[2]);
and and4(OUT[3], A[3] , B[3]);
and and5(OUT[4], A[4] , B[4]);
and and6(OUT[5], A[5] , B[5]);
and and7(OUT[6], A[6] , B[6]);
and and8(OUT[7], A[7] , B[7]);
and and9(OUT[8], A[8] , B[8]);
and and10(OUT[9], A[9] , B[9]);
and and11(OUT[10], A[10] , B[10]);
and and12(OUT[11], A[11] , B[11]);
and and13(OUT[12], A[12] , B[12]);
and and14(OUT[13], A[13] , B[13]);
and and15(OUT[14], A[14] , B[14]);
and and16(OUT[15], A[15] , B[15]);
and and17(OUT[16], A[16] , B[16]);
and and18(OUT[17], A[17] , B[17]);
and and19(OUT[18], A[18] , B[18]);
and and20(OUT[19], A[19] , B[19]);
and and21(OUT[20], A[20] , B[20]);
and and22(OUT[21], A[21] , B[21]);
and and23(OUT[22], A[22] , B[22]);
and and24(OUT[23], A[23] , B[23]);
and and25(OUT[24], A[24] , B[24]);
and and26(OUT[25], A[25] , B[25]);
and and27(OUT[26], A[26] , B[26]);
and and28(OUT[27], A[27] , B[27]);
and and29(OUT[28], A[28] , B[28]);
and and30(OUT[29], A[29] , B[29]);
and and31(OUT[30], A[30] , B[30]);
and and32(OUT[31], A[31] , B[31]);


endmodule