library verilog;
use verilog.vl_types.all;
entity set_less_than_32_testbench is
end set_less_than_32_testbench;
