library verilog;
use verilog.vl_types.all;
entity mux_4x1_testbench is
end mux_4x1_testbench;
