library verilog;
use verilog.vl_types.all;
entity adder_1_bit_testbench is
end adder_1_bit_testbench;
