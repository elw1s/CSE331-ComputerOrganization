library verilog;
use verilog.vl_types.all;
entity and_32_bit_testbench is
end and_32_bit_testbench;
