
module not_32_bit(input [31:0] A , output[31:0] OUT);



not F1(OUT[0] , A[0]);
not F2(OUT[1] , A[1]);
not F3(OUT[2] , A[2]);
not F4(OUT[3] , A[3]);
not F5(OUT[4] , A[4]);
not F6(OUT[5] , A[5]);
not F7(OUT[6] , A[6]);
not F8(OUT[7] , A[7]);
not F9(OUT[8] , A[8]);
not F10(OUT[9] , A[9]);
not F11(OUT[10] , A[10]);
not F12(OUT[11] , A[11]);
not F13(OUT[12] , A[12]);
not F14(OUT[13] , A[13]);
not F15(OUT[14] , A[14]);
not F16(OUT[15] , A[15]);
not F17(OUT[16] , A[16]);
not F18(OUT[17] , A[17]);
not F19(OUT[18] , A[18]);
not F20(OUT[19] , A[19]);
not F21(OUT[20] , A[20]);
not F22(OUT[21] , A[21]);
not F23(OUT[22] , A[22]);
not F24(OUT[23] , A[23]);
not F25(OUT[24] , A[24]);
not F26(OUT[25] , A[25]);
not F27(OUT[26] , A[26]);
not F28(OUT[27] , A[27]);
not F29(OUT[28] , A[28]);
not F30(OUT[29] , A[29]);
not F31(OUT[30] , A[30]);
not F32(OUT[31] , A[31]);

endmodule