library verilog;
use verilog.vl_types.all;
entity xor_32_bit_testbench is
end xor_32_bit_testbench;
