library verilog;
use verilog.vl_types.all;
entity or_32_bit_testbench is
end or_32_bit_testbench;
