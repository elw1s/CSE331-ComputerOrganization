library verilog;
use verilog.vl_types.all;
entity nor_32_bit_testbench is
end nor_32_bit_testbench;
