library verilog;
use verilog.vl_types.all;
entity mux_8x1_testbench is
end mux_8x1_testbench;
