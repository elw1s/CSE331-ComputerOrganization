library verilog;
use verilog.vl_types.all;
entity and_6bit is
    port(
        A               : in     vl_logic;
        B               : in     vl_logic;
        C               : in     vl_logic;
        D               : in     vl_logic;
        E               : in     vl_logic;
        F               : in     vl_logic;
        \OUT\           : out    vl_logic
    );
end and_6bit;
