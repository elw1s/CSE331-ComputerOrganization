library verilog;
use verilog.vl_types.all;
entity mux_2x1_testbench is
end mux_2x1_testbench;
