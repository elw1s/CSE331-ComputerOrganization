library verilog;
use verilog.vl_types.all;
entity ProgramCounterTestBench is
end ProgramCounterTestBench;
