library verilog;
use verilog.vl_types.all;
entity instruction_memory_testbench is
end instruction_memory_testbench;
