library verilog;
use verilog.vl_types.all;
entity mips_16bit_testbench is
end mips_16bit_testbench;
