library verilog;
use verilog.vl_types.all;
entity adder_32_bit_testbench is
end adder_32_bit_testbench;
