library verilog;
use verilog.vl_types.all;
entity control_testbench is
end control_testbench;
