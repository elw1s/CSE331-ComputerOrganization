library verilog;
use verilog.vl_types.all;
entity xorgate_testbench is
end xorgate_testbench;
