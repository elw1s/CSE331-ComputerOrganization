library verilog;
use verilog.vl_types.all;
entity mux_8x1_32bit_testbench is
end mux_8x1_32bit_testbench;
